library ieee;
use ieee.std_logic_1164.all;

package Ram_Pkg is
    type RamVector is array (0 to 255) of std_logic_vector(7 downto 0);
end Ram_Pkg;

package body Ram_Pkg is
end Ram_Pkg;
